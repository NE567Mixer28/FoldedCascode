** sch_path: /home/ttuser/FoldedCascode_OTA/xschem/OTA_FoldedCascode_L.sch
.subckt OTA_FoldedCascode_L IN+ IN- OUT VDD GND Vc Vp
*.PININFO IN+:I IN-:I OUT:O VDD:B GND:B Vc:B Vp:B
XM1 D1 IN+ S S sky130_fd_pr__pfet_01v8 L=1 W=10 nf=1 m=5
XM2 D2 IN- S S sky130_fd_pr__pfet_01v8 L=1 W=10 nf=1 m=5
XM3 D1 Vc GND GND sky130_fd_pr__nfet_01v8 L=10 W=2 nf=1 m=1
XM4 D2 Vc GND GND sky130_fd_pr__nfet_01v8 L=10 W=2 nf=1 m=1
XM5 G Vc D1 GND sky130_fd_pr__nfet_01v8 L=2 W=3 nf=1 m=1
XM6 OUT Vc D2 GND sky130_fd_pr__nfet_01v8 L=2 W=3 nf=1 m=1
XM7 G Vc D9 D9 sky130_fd_pr__pfet_01v8 L=5 W=10 nf=1 m=1
XM8 OUT Vc D10 D10 sky130_fd_pr__pfet_01v8 L=5 W=10 nf=1 m=1
XM9 D9 G VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=26 nf=1 m=1
XM10 D10 G VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=26 nf=1 m=1
XM11 S Vp net1 VDD sky130_fd_pr__pfet_01v8 L=5 W=5 nf=1 m=1
XM12 net1 Vp VDD VDD sky130_fd_pr__pfet_01v8 L=5 W=5 nf=1 m=1
XR5 GND Vc GND sky130_fd_pr__res_xhigh_po W=0.35 L=3.2 mult=1 m=1
XR1 Vc VDD GND sky130_fd_pr__res_xhigh_po W=0.35 L=5 mult=1 m=1
XR2 Vp VDD GND sky130_fd_pr__res_xhigh_po W=0.35 L=5 mult=1 m=1
XR3 GND Vp GND sky130_fd_pr__res_xhigh_po W=0.35 L=1.94 mult=1 m=1
.ends
.end
